----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:56:41 04/24/2019 
-- Design Name: 
-- Module Name:    the_other_mem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
----------------------- ENTITY --------------------------------------------
entity memory is
	port
	(
		address: in std_logic_vector (31 downto 0); --ADDRESS TO WRITE OR READ
		data_write: in std_logic_vector (31 downto 0); -- DATA TO BE WRITTEN
		memWrite: in std_logic; --HIGH FOR WRITING 
		memRead: in std_logic; --HIGH FOR READING
		--clk: in std_logic; -- CLOCK
		data_read: out std_logic_vector (31 downto 0) --DATA FROM ADDRESS address
	);
end memory;

architecture memory1 of memory is
	
	--TYPE of memory section
	type MEMORY_ARRAY is array (0 to 31) of std_logic_vector (31 downto 0);
	
	-- MEMORY
	signal data: MEMORY_ARRAY := (
X"00221820",
X"8D010000",	--LW reg1, offset (0); reg1 = 0, offset 0
X"00000000", 
X"00000000",
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000", 
X"00000000", 
X"00000000",
X"00000000",
X"00000000");


	signal fakeaddress: std_logic_vector(31 downto 0):= (others => '0');
	--GENERAL CONSTANTS
	constant CONST_ZERO: std_logic_vector(31 downto 0):= (others => '0');
		
	
	begin
		process (address, memRead, data_write) 
		begin
				if( address(0) /= '0' and address(0) /= '1')then
					data_read <= CONST_ZERO;
				elsif(memRead = '1' AND memWrite = '1') then -- if both memREAD and memWRITE are ON, there is a problem, so I put 0 in OUTPUT
					data_read <= CONST_ZERO;
				elsif( memRead = '1') then	 --if I want to read data										
					data_read <= data( conv_integer( unsigned( address ) )/4 );
				elsif (memWrite = '1') then -- if I want to write data					
					data( conv_integer( unsigned( address ) )/4 )<= data_write;
			
				end if;

		end process;
	
end memory1;